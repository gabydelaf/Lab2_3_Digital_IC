Library IEEE;
use IEEE.std_logic_1164.all;

Entity signal_mapper is 
  Port (sseg_out : In std_logic(6 downto 0);
        a, b, c, d, e, f, g : Out std_logic);
End signal_mapper;

Architecture of signal_mapper Is
  a <= sseg_out(0);
  b <= sseg_out(1);
  c <= sseg_out(2);
  d <= sseg_out(3);
  e <= sseg_out(4);
  f <= sseg_out(5);
  g <= sseg_out(6);
End Architecture signal_mapper;
